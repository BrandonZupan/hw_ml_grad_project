// multiply.v

module multiply (
    input [255:0]   op0_value;
    input [255:0]   op1_value;

    input [2:0]     vlmul;

    output [255:0]  mul_out;
);

endmodule